`timescale 1ns / 1ps

module hello;
    initial begin
        $display("🚀 Hello, Verilog! Starting my 15-day challenge.");
        $finish;
    end
endmodule
